module inv(A,Z);
  input A;
  output Z;

  assign Z = ~A;
endmodule
